package fifo_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"
   

  `include "fifo_trans.sv"
  `include "fifo_driver.sv"
  `include "fifo_monitor.sv"
  `include "fifo_seqr.sv"
  `include "fifo_base_seqs.sv"
  `include "fifo_agent.sv"
  `include "fifo_scoreboard.sv"
  
 `include "fifo_virtual_seqr.sv"
  `include "fifo_base_vseqs.sv" 
   
  
 `include "fifo_env.sv"
  
 `include "fifo_base_test.sv"
  
 //reset test
 `include "fifo_reset_seqs.sv"
 `include "fifo_reset_vseqs.sv"
 `include "fifo_reset_test.sv"

 //overflow test
  `include "fifo_buf_full_seqs.sv"
  `include "fifo_full_vseqs.sv"
  `include "fifo_full_test.sv"
  

  
endpackage
